library ieee;
USE ieee.std_logic_1164.ALL;

package myPackages is
  type Block_Cache is array (7 downto 0) of std_logic_vector(15 downto 0);
  type Cache is array (31 downto 0) of Block_Cache;
  type Taglist is array (31 downto 0) of std_logic_vector(2 downto 0);
end package;

library ieee;
USE ieee.std_logic_1164.ALL;
--use IEEE.std_logic_arith.all;
use ieee.numeric_std.all;

use work.myPackages.all;

Entity Cache_DataMemory is
	PORT (clk : IN std_logic;
	      MR, MW, RamRead, NoWrite,rst,int : IN std_logic;
	      add : IN std_logic_vector(7 DOWNTO 0);
	      datain : IN std_logic_vector(31 DOWNTO 0);
	      dataout : OUT std_logic_vector(31 DOWNTO 0);
	      blockIN: IN Block_Cache;
	      blockOUT: OUT Block_Cache);
END Cache_DataMemory;

ARCHITECTURE combinational OF Cache_DataMemory IS

SIGNAL storage : Cache;
signal address: std_logic_vector(7 DOWNTO 0);
Begin
process(rst,int,add)
begin
if rst = '1' then 
address <= "00000000";
elsif int = '1' then 
address <= "00000010";
else
address <= add;
end if;
end process;
blockOUT<= storage(to_integer(unsigned(address(7 downto 3))));
process(clk)
	variable index, displacement: Integer;
	begin
	index:= to_integer(unsigned(address(7 downto 3)));
	displacement:= to_integer(unsigned(address(2 downto 0)));
	IF falling_edge(clk) then 
		if MW = '1' and NoWrite = '0' and RamRead = '0' THEN  
		storage(index)(displacement)<= datain(15 downto 0); storage(index)(displacement+1)<= datain(31 downto 16);
		elsif  RamRead = '1' then 
		storage(index) <= blockIN;
		end if;
	END IF;
END PROCESS;

process(MR, storage, address)
	variable index, displacement: Integer;
	begin
	index:= to_integer(unsigned(address(7 downto 3)));
	displacement:= to_integer(unsigned(address(2 downto 0)));
	if MR = '1' or rst='1' or int='1' then dataout <= storage(index)(displacement+1)&storage(index)(displacement);
	else dataout <=(others=>'0');
	end if;
end process;

End ARCHITECTURE;

library ieee;
USE ieee.std_logic_1164.ALL;
--use IEEE.std_logic_arith.all;
use ieee.numeric_std.all;

use work.myPackages.all;

Entity Cache_InstructionMemory is
	PORT (clk : IN std_logic;
	      MW, RamRead, nowrite: IN std_logic;
	      address, addressWrite : IN std_logic_vector(7 DOWNTO 0);
	      datain : IN std_logic_vector (1 DOWNTO 0);
	      dataout : OUT std_logic_vector(15 DOWNTO 0);
	      blockIN: IN Block_Cache
	      );
END Cache_InstructionMemory;

ARCHITECTURE combinational2 OF Cache_InstructionMemory IS

SIGNAL storage : Cache;
Begin

process(clk)
	variable index, displacement, indexread: Integer;
	begin
	index:= to_integer(unsigned(addressWrite(7 downto 3)));
	displacement:=to_integer(unsigned(addressWrite(2 downto 0)));
	indexread:= to_integer(unsigned(address(7 downto 3)));
	IF falling_edge(clk) then 
		if MW = '1' and NoWrite = '0' and RamRead = '0' THEN  
		storage(index)(displacement)(15 downto 14)<= datain;
		elsif  RamRead = '1' then 
		storage(indexread) <= blockIN;
		end if;
	END IF;
END PROCESS;

process(storage, address)
	variable index, displacement: Integer;
	begin
	index:= to_integer(unsigned(address(7 downto 3)));
	displacement:= to_integer(unsigned(address(2 downto 0)));
	dataout <= storage(index)(displacement);
end process;

End ARCHITECTURE;

library ieee;
USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;

use work.myPackages.all;

Entity Cache_Controller is
	PORT (clk, Vrst, rst, MR, MW, MWInstr,int: IN std_logic;
	      add, addressInstr, addressInstrWrite : IN std_logic_vector(10 DOWNTO 3);
	      AddressToRam: OUT std_logic_vector(10 DOWNTO 0);
	      MemW, CacheW, CacheWInstr, ignore: OUT std_logic);
END Cache_Controller;

ARCHITECTURE control OF Cache_Controller IS

signal TagArray, TagArrinstr : Taglist;
signal ValidArray, dirtyArray, ValidArrInstr : std_logic_vector(31 downto 0);
signal TagWrite, dirtyWrite, TagWriteInstr: std_logic;
signal index, indexInstr, indexInstrWrite: Integer;
signal tag,tagInstr, tagInstrWrite : std_logic_vector(2 downto 0);
signal address: std_logic_vector(10 downto 3);
Begin
tag<= address(10 downto 8);
tagInstr<= addressInstr(10 downto 8);
tagInstrWrite<= addressInstrWrite(10 downto 8);
index<= to_integer(unsigned((address(7 downto 3))));
indexInstr<= to_integer(unsigned((addressInstr(7 downto 3))));
indexInstrWrite<= to_integer(unsigned((addressInstrWrite(7 downto 3))));
process(rst,int,add)
begin
if rst = '1' then 
address <= "00000000";
elsif int = '1' then 
address <= "00000010";
else
address <= add;
end if;
end process;
process(clk,MR, MW, address, TagArray, ValidArray, dirtyArray, rst, ValidArrInstr, TagArrinstr,addressInstr,addressInstrWrite,MWInstr)
variable dataMissPrior: integer;
begin

dataMissPrior:=0;
--CacheW<='0'; TagWrite<='0';
if rising_edge(clk) then
	MemW<='0'; CacheW<='0'; TagWrite<='0'; dirtyWrite <= '0'; CacheWInstr <='0'; TagWriteInstr<='0'; ignore<='0';
	if MR ='1' or MW = '1' or rst='1' or int='1' then 
		   if (ValidArray(index) = '0' or TagArray(index) /= tag) then   dataMissPrior :=1;   -- Miss
			if dirtyArray(index) = '0' then  CacheW<= '1'; TagWrite<='1'; AddressToRam<=address(10 downto 3)&"000";
			else MemW<= '1'; dirtyWrite<= '1'; AddressToRam<=TagArray(index)&Address(7 downto 3)&"000";
			end if;
		   end if;
	end if;
		
	if dataMissPrior = 0 then
		if (ValidArrInstr(indexInstr) = '0' or TagArrinstr(indexInstr) /= tagInstr) and addressInstr /= "UUUUUUUU" and addressInstr /= "XXXXXXXX" then 
				CacheWInstr <='1'; TagWriteInstr<='1'; AddressToRam<=addressInstr(10 downto 3)&"000"; end if;
		if MWInstr ='1' and (ValidArrInstr(indexInstrWrite) = '0' or TagArrinstr(indexInstrWrite) /= tagInstrWrite) then
			ignore <='1';
		end if;
			
	end if;
	
end if;
end process;

process (clk, rst, tagWrite, address, dirtyWrite, addressInstr,TagWriteInstr)
	begin
	if Vrst ='1' then  ValidArray<=(others=>'0'); dirtyArray<=(others=>'0'); ValidArrInstr<=(others=>'0'); end if;
	if falling_edge(clk) then 
		if dirtyWrite = '1' then dirtyArray(index)<= '0'; end if; 
 
		if MW = '1' and ValidArray(index) = '1' and TagArray(index) = tag then -- Write HIT
			dirtyArray(index)<= '1'; end if;
		if tagWrite = '1' then TagArray(index) <= tag; ValidArray(index)<='1'; end if;
		if TagWriteInstr ='1' then TagArrinstr(indexInstr) <=tagInstr; ValidArrInstr(indexInstr)<='1'; end if;
	end if;
end process;

End control;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;
use work.myPackages.all;

ENTITY MainMemory IS

PORT (clk, we : IN std_logic;
address : IN std_logic_vector(10 DOWNTO 0);
datain : IN Block_Cache;
dataout : OUT Block_Cache);
END MainMemory;

ARCHITECTURE main OF MainMemory IS

TYPE ram_type IS ARRAY(0 TO 2047) of std_logic_vector(15 DOWNTO 0);

SIGNAL ram : ram_type := (
0=> "0000000000010000" ,
1=> "0000000000000000" ,
2=> "0000000100000000" ,
3=> "0000000000000000" ,
4=> "0011100000000000" ,
5=> "0000000100000000" ,
6=> "0011110000000000" ,
7=> "0000000000000010" ,
8=> "0001000000000000" ,
9=> "0001000000000000" ,
10=> "0001000000000000" ,
11=> "0001000000000000" ,
12=> "0001000000000000" ,
13=> "0001000000000000" ,
14=> "0001000000000000" ,
15=> "0001000000000000" ,
16=> "0001101001000001" ,
17=> "0001101010000010" ,
18=> "0001101011000011" ,
19=> "0001101100000100" ,
20=> "0001101110000110" ,
21=> "0001101111000111" ,
22=> "0011000100000000" ,
23=> "0010001001000000" ,
24=> "0001010111000111" ,
25=> "0001000000000000" ,
26=> "0001000000000000" ,
27=> "0001000000000000" ,
28=> "0001000000000000" ,
29=> "0001000000000000" ,
30=> "0001000000000000" ,
31=> "0001000000000000" ,
32=> "0001000000000000" ,
33=> "0001000000000000" ,
34=> "0001000000000000" ,
35=> "0001000000000000" ,
36=> "0001000000000000" ,
37=> "0001000000000000" ,
38=> "0001000000000000" ,
39=> "0001000000000000" ,
40=> "0001000000000000" ,
41=> "0001000000000000" ,
42=> "0001000000000000" ,
43=> "0001000000000000" ,
44=> "0001000000000000" ,
45=> "0001000000000000" ,
46=> "0001000000000000" ,
47=> "0001000000000000" ,
48=> "0000100001101101" ,
49=> "0010000010000000" ,
50=> "0001010111000111" ,
51=> "0001000000000000" ,
52=> "0001000000000000" ,
53=> "0001000000000000" ,
54=> "0001000000000000" ,
55=> "0001000000000000" ,
56=> "0001000000000000" ,
57=> "0001000000000000" ,
58=> "0001000000000000" ,
59=> "0001000000000000" ,
60=> "0001000000000000" ,
61=> "0001000000000000" ,
62=> "0001000000000000" ,
63=> "0001000000000000" ,
64=> "0001000000000000" ,
65=> "0001000000000000" ,
66=> "0001000000000000" ,
67=> "0001000000000000" ,
68=> "0001000000000000" ,
69=> "0001000000000000" ,
70=> "0001000000000000" ,
71=> "0001000000000000" ,
72=> "0001000000000000" ,
73=> "0001000000000000" ,
74=> "0001000000000000" ,
75=> "0001000000000000" ,
76=> "0001000000000000" ,
77=> "0001000000000000" ,
78=> "0001000000000000" ,
79=> "0001000000000000" ,
80=> "0010000011000000" ,
81=> "0001001101000101" ,
82=> "0001010101000101" ,
83=> "0001101110000110" ,
84=> "0010000110000000" ,
85=> "0001010001000001" ,
86=> "0001000000000000" ,
87=> "0001000000000000" ,
88=> "0001000000000000" ,
89=> "0001000000000000" ,
90=> "0001000000000000" ,
91=> "0001000000000000" ,
92=> "0001000000000000" ,
93=> "0001000000000000" ,
94=> "0001000000000000" ,
95=> "0001000000000000" ,
96=> "0001000000000000" ,
97=> "0001000000000000" ,
98=> "0001000000000000" ,
99=> "0001000000000000" ,
100=> "0001000000000000" ,
101=> "0001000000000000" ,
102=> "0001000000000000" ,
103=> "0001000000000000" ,
104=> "0001000000000000" ,
105=> "0001000000000000" ,
106=> "0001000000000000" ,
107=> "0001000000000000" ,
108=> "0001000000000000" ,
109=> "0001000000000000" ,
110=> "0001000000000000" ,
111=> "0001000000000000" ,
112=> "0001000000000000" ,
113=> "0001000000000000" ,
114=> "0001000000000000" ,
115=> "0001000000000000" ,
116=> "0001000000000000" ,
117=> "0001000000000000" ,
118=> "0001000000000000" ,
119=> "0001000000000000" ,
120=> "0001000000000000" ,
121=> "0001000000000000" ,
122=> "0001000000000000" ,
123=> "0001000000000000" ,
124=> "0001000000000000" ,
125=> "0001000000000000" ,
126=> "0001000000000000" ,
127=> "0001000000000000" ,
128=> "0001000000000000" ,
129=> "0001000000000000" ,
130=> "0001000000000000" ,
131=> "0001000000000000" ,
132=> "0001000000000000" ,
133=> "0001000000000000" ,
134=> "0001000000000000" ,
135=> "0001000000000000" ,
136=> "0001000000000000" ,
137=> "0001000000000000" ,
138=> "0001000000000000" ,
139=> "0001000000000000" ,
140=> "0001000000000000" ,
141=> "0001000000000000" ,
142=> "0001000000000000" ,
143=> "0001000000000000" ,
144=> "0001000000000000" ,
145=> "0001000000000000" ,
146=> "0001000000000000" ,
147=> "0001000000000000" ,
148=> "0001000000000000" ,
149=> "0001000000000000" ,
150=> "0001000000000000" ,
151=> "0001000000000000" ,
152=> "0001000000000000" ,
153=> "0001000000000000" ,
154=> "0001000000000000" ,
155=> "0001000000000000" ,
156=> "0001000000000000" ,
157=> "0001000000000000" ,
158=> "0001000000000000" ,
159=> "0001000000000000" ,
160=> "0001000000000000" ,
161=> "0001000000000000" ,
162=> "0001000000000000" ,
163=> "0001000000000000" ,
164=> "0001000000000000" ,
165=> "0001000000000000" ,
166=> "0001000000000000" ,
167=> "0001000000000000" ,
168=> "0001000000000000" ,
169=> "0001000000000000" ,
170=> "0001000000000000" ,
171=> "0001000000000000" ,
172=> "0001000000000000" ,
173=> "0001000000000000" ,
174=> "0001000000000000" ,
175=> "0001000000000000" ,
176=> "0001000000000000" ,
177=> "0001000000000000" ,
178=> "0001000000000000" ,
179=> "0001000000000000" ,
180=> "0001000000000000" ,
181=> "0001000000000000" ,
182=> "0001000000000000" ,
183=> "0001000000000000" ,
184=> "0001000000000000" ,
185=> "0001000000000000" ,
186=> "0001000000000000" ,
187=> "0001000000000000" ,
188=> "0001000000000000" ,
189=> "0001000000000000" ,
190=> "0001000000000000" ,
191=> "0001000000000000" ,
192=> "0001000000000000" ,
193=> "0001000000000000" ,
194=> "0001000000000000" ,
195=> "0001000000000000" ,
196=> "0001000000000000" ,
197=> "0001000000000000" ,
198=> "0001000000000000" ,
199=> "0001000000000000" ,
200=> "0001000000000000" ,
201=> "0001000000000000" ,
202=> "0001000000000000" ,
203=> "0001000000000000" ,
204=> "0001000000000000" ,
205=> "0001000000000000" ,
206=> "0001000000000000" ,
207=> "0001000000000000" ,
208=> "0001000000000000" ,
209=> "0001000000000000" ,
210=> "0001000000000000" ,
211=> "0001000000000000" ,
212=> "0001000000000000" ,
213=> "0001000000000000" ,
214=> "0001000000000000" ,
215=> "0001000000000000" ,
216=> "0001000000000000" ,
217=> "0001000000000000" ,
218=> "0001000000000000" ,
219=> "0001000000000000" ,
220=> "0001000000000000" ,
221=> "0001000000000000" ,
222=> "0001000000000000" ,
223=> "0001000000000000" ,
224=> "0001000000000000" ,
225=> "0001000000000000" ,
226=> "0001000000000000" ,
227=> "0001000000000000" ,
228=> "0001000000000000" ,
229=> "0001000000000000" ,
230=> "0001000000000000" ,
231=> "0001000000000000" ,
232=> "0001000000000000" ,
233=> "0001000000000000" ,
234=> "0001000000000000" ,
235=> "0001000000000000" ,
236=> "0001000000000000" ,
237=> "0001000000000000" ,
238=> "0001000000000000" ,
239=> "0001000000000000" ,
240=> "0001000000000000" ,
241=> "0001000000000000" ,
242=> "0001000000000000" ,
243=> "0001000000000000" ,
244=> "0001000000000000" ,
245=> "0001000000000000" ,
246=> "0001000000000000" ,
247=> "0001000000000000" ,
248=> "0001000000000000" ,
249=> "0001000000000000" ,
250=> "0001000000000000" ,
251=> "0001000000000000" ,
252=> "0001000000000000" ,
253=> "0001000000000000" ,
254=> "0001000000000000" ,
255=> "0001000000000000" ,
256=> "0000001000000000" ,
257=> "0001100110000110" ,
258=> "0010101000000000" ,
259=> "0001000000000000" ,
260=> "0001000000000000" ,
261=> "0001000000000000" ,
262=> "0001000000000000" ,
263=> "0001000000000000" ,
264=> "0001000000000000" ,
265=> "0001000000000000" ,
266=> "0001000000000000" ,
267=> "0001000000000000" ,
268=> "0001000000000000" ,
269=> "0001000000000000" ,
270=> "0001000000000000" ,
271=> "0001000000000000" ,
272=> "0001000000000000" ,
273=> "0001000000000000" ,
274=> "0001000000000000" ,
275=> "0001000000000000" ,
276=> "0001000000000000" ,
277=> "0001000000000000" ,
278=> "0001000000000000" ,
279=> "0001000000000000" ,
280=> "0001000000000000" ,
281=> "0001000000000000" ,
282=> "0001000000000000" ,
283=> "0001000000000000" ,
284=> "0001000000000000" ,
285=> "0001000000000000" ,
286=> "0001000000000000" ,
287=> "0001000000000000" ,
288=> "0001000000000000" ,
289=> "0001000000000000" ,
290=> "0001000000000000" ,
291=> "0001000000000000" ,
292=> "0001000000000000" ,
293=> "0001000000000000" ,
294=> "0001000000000000" ,
295=> "0001000000000000" ,
296=> "0001000000000000" ,
297=> "0001000000000000" ,
298=> "0001000000000000" ,
299=> "0001000000000000" ,
300=> "0001000000000000" ,
301=> "0001000000000000" ,
302=> "0001000000000000" ,
303=> "0001000000000000" ,
304=> "0001000000000000" ,
305=> "0001000000000000" ,
306=> "0001000000000000" ,
307=> "0001000000000000" ,
308=> "0001000000000000" ,
309=> "0001000000000000" ,
310=> "0001000000000000" ,
311=> "0001000000000000" ,
312=> "0001000000000000" ,
313=> "0001000000000000" ,
314=> "0001000000000000" ,
315=> "0001000000000000" ,
316=> "0001000000000000" ,
317=> "0001000000000000" ,
318=> "0001000000000000" ,
319=> "0001000000000000" ,
320=> "0001000000000000" ,
321=> "0001000000000000" ,
322=> "0001000000000000" ,
323=> "0001000000000000" ,
324=> "0001000000000000" ,
325=> "0001000000000000" ,
326=> "0001000000000000" ,
327=> "0001000000000000" ,
328=> "0001000000000000" ,
329=> "0001000000000000" ,
330=> "0001000000000000" ,
331=> "0001000000000000" ,
332=> "0001000000000000" ,
333=> "0001000000000000" ,
334=> "0001000000000000" ,
335=> "0001000000000000" ,
336=> "0001000000000000" ,
337=> "0001000000000000" ,
338=> "0001000000000000" ,
339=> "0001000000000000" ,
340=> "0001000000000000" ,
341=> "0001000000000000" ,
342=> "0001000000000000" ,
343=> "0001000000000000" ,
344=> "0001000000000000" ,
345=> "0001000000000000" ,
346=> "0001000000000000" ,
347=> "0001000000000000" ,
348=> "0001000000000000" ,
349=> "0001000000000000" ,
350=> "0001000000000000" ,
351=> "0001000000000000" ,
352=> "0001000000000000" ,
353=> "0001000000000000" ,
354=> "0001000000000000" ,
355=> "0001000000000000" ,
356=> "0001000000000000" ,
357=> "0001000000000000" ,
358=> "0001000000000000" ,
359=> "0001000000000000" ,
360=> "0001000000000000" ,
361=> "0001000000000000" ,
362=> "0001000000000000" ,
363=> "0001000000000000" ,
364=> "0001000000000000" ,
365=> "0001000000000000" ,
366=> "0001000000000000" ,
367=> "0001000000000000" ,
368=> "0001000000000000" ,
369=> "0001000000000000" ,
370=> "0001000000000000" ,
371=> "0001000000000000" ,
372=> "0001000000000000" ,
373=> "0001000000000000" ,
374=> "0001000000000000" ,
375=> "0001000000000000" ,
376=> "0001000000000000" ,
377=> "0001000000000000" ,
378=> "0001000000000000" ,
379=> "0001000000000000" ,
380=> "0001000000000000" ,
381=> "0001000000000000" ,
382=> "0001000000000000" ,
383=> "0001000000000000" ,
384=> "0001000000000000" ,
385=> "0001000000000000" ,
386=> "0001000000000000" ,
387=> "0001000000000000" ,
388=> "0001000000000000" ,
389=> "0001000000000000" ,
390=> "0001000000000000" ,
391=> "0001000000000000" ,
392=> "0001000000000000" ,
393=> "0001000000000000" ,
394=> "0001000000000000" ,
395=> "0001000000000000" ,
396=> "0001000000000000" ,
397=> "0001000000000000" ,
398=> "0001000000000000" ,
399=> "0001000000000000" ,
400=> "0001000000000000" ,
401=> "0001000000000000" ,
402=> "0001000000000000" ,
403=> "0001000000000000" ,
404=> "0001000000000000" ,
405=> "0001000000000000" ,
406=> "0001000000000000" ,
407=> "0001000000000000" ,
408=> "0001000000000000" ,
409=> "0001000000000000" ,
410=> "0001000000000000" ,
411=> "0001000000000000" ,
412=> "0001000000000000" ,
413=> "0001000000000000" ,
414=> "0001000000000000" ,
415=> "0001000000000000" ,
416=> "0001000000000000" ,
417=> "0001000000000000" ,
418=> "0001000000000000" ,
419=> "0001000000000000" ,
420=> "0001000000000000" ,
421=> "0001000000000000" ,
422=> "0001000000000000" ,
423=> "0001000000000000" ,
424=> "0001000000000000" ,
425=> "0001000000000000" ,
426=> "0001000000000000" ,
427=> "0001000000000000" ,
428=> "0001000000000000" ,
429=> "0001000000000000" ,
430=> "0001000000000000" ,
431=> "0001000000000000" ,
432=> "0001000000000000" ,
433=> "0001000000000000" ,
434=> "0001000000000000" ,
435=> "0001000000000000" ,
436=> "0001000000000000" ,
437=> "0001000000000000" ,
438=> "0001000000000000" ,
439=> "0001000000000000" ,
440=> "0001000000000000" ,
441=> "0001000000000000" ,
442=> "0001000000000000" ,
443=> "0001000000000000" ,
444=> "0001000000000000" ,
445=> "0001000000000000" ,
446=> "0001000000000000" ,
447=> "0001000000000000" ,
448=> "0001000000000000" ,
449=> "0001000000000000" ,
450=> "0001000000000000" ,
451=> "0001000000000000" ,
452=> "0001000000000000" ,
453=> "0001000000000000" ,
454=> "0001000000000000" ,
455=> "0001000000000000" ,
456=> "0001000000000000" ,
457=> "0001000000000000" ,
458=> "0001000000000000" ,
459=> "0001000000000000" ,
460=> "0001000000000000" ,
461=> "0001000000000000" ,
462=> "0001000000000000" ,
463=> "0001000000000000" ,
464=> "0001000000000000" ,
465=> "0001000000000000" ,
466=> "0001000000000000" ,
467=> "0001000000000000" ,
468=> "0001000000000000" ,
469=> "0001000000000000" ,
470=> "0001000000000000" ,
471=> "0001000000000000" ,
472=> "0001000000000000" ,
473=> "0001000000000000" ,
474=> "0001000000000000" ,
475=> "0001000000000000" ,
476=> "0001000000000000" ,
477=> "0001000000000000" ,
478=> "0001000000000000" ,
479=> "0001000000000000" ,
480=> "0001000000000000" ,
481=> "0001000000000000" ,
482=> "0001000000000000" ,
483=> "0001000000000000" ,
484=> "0001000000000000" ,
485=> "0001000000000000" ,
486=> "0001000000000000" ,
487=> "0001000000000000" ,
488=> "0001000000000000" ,
489=> "0001000000000000" ,
490=> "0001000000000000" ,
491=> "0001000000000000" ,
492=> "0001000000000000" ,
493=> "0001000000000000" ,
494=> "0001000000000000" ,
495=> "0001000000000000" ,
496=> "0001000000000000" ,
497=> "0001000000000000" ,
498=> "0001000000000000" ,
499=> "0001000000000000" ,
500=> "0001000000000000" ,
501=> "0001000000000000" ,
502=> "0001000000000000" ,
503=> "0001000000000000" ,
504=> "0001000000000000" ,
505=> "0001000000000000" ,
506=> "0001000000000000" ,
507=> "0001000000000000" ,
508=> "0001000000000000" ,
509=> "0001000000000000" ,
510=> "0001000000000000" ,
511=> "0001000000000000" ,
512=> "0011001000000110" ,
513=> "0010010110000000" ,
514=> "0001010110000110" ,
515=> "0001000000000000" ,
516=> "0001000000000000" ,
517=> "0001000000000000" ,
518=> "0001000000000000" ,
519=> "0001000000000000" ,
520=> "0001000000000000" ,
521=> "0001000000000000" ,
522=> "0001000000000000" ,
523=> "0001000000000000" ,
524=> "0001000000000000" ,
525=> "0001000000000000" ,
526=> "0001000000000000" ,
527=> "0001000000000000" ,
528=> "0001000000000000" ,
529=> "0001000000000000" ,
530=> "0001000000000000" ,
531=> "0001000000000000" ,
532=> "0001000000000000" ,
533=> "0001000000000000" ,
534=> "0001000000000000" ,
535=> "0001000000000000" ,
536=> "0001000000000000" ,
537=> "0001000000000000" ,
538=> "0001000000000000" ,
539=> "0001000000000000" ,
540=> "0001000000000000" ,
541=> "0001000000000000" ,
542=> "0001000000000000" ,
543=> "0001000000000000" ,
544=> "0001000000000000" ,
545=> "0001000000000000" ,
546=> "0001000000000000" ,
547=> "0001000000000000" ,
548=> "0001000000000000" ,
549=> "0001000000000000" ,
550=> "0001000000000000" ,
551=> "0001000000000000" ,
552=> "0001000000000000" ,
553=> "0001000000000000" ,
554=> "0001000000000000" ,
555=> "0001000000000000" ,
556=> "0001000000000000" ,
557=> "0001000000000000" ,
558=> "0001000000000000" ,
559=> "0001000000000000" ,
560=> "0001000000000000" ,
561=> "0001000000000000" ,
562=> "0001000000000000" ,
563=> "0001000000000000" ,
564=> "0001000000000000" ,
565=> "0001000000000000" ,
566=> "0001000000000000" ,
567=> "0001000000000000" ,
568=> "0001000000000000" ,
569=> "0001000000000000" ,
570=> "0001000000000000" ,
571=> "0001000000000000" ,
572=> "0001000000000000" ,
573=> "0001000000000000" ,
574=> "0001000000000000" ,
575=> "0001000000000000" ,
576=> "0001000000000000" ,
577=> "0001000000000000" ,
578=> "0001000000000000" ,
579=> "0001000000000000" ,
580=> "0001000000000000" ,
581=> "0001000000000000" ,
582=> "0001000000000000" ,
583=> "0001000000000000" ,
584=> "0001000000000000" ,
585=> "0001000000000000" ,
586=> "0001000000000000" ,
587=> "0001000000000000" ,
588=> "0001000000000000" ,
589=> "0001000000000000" ,
590=> "0001000000000000" ,
591=> "0001000000000000" ,
592=> "0001000000000000" ,
593=> "0001000000000000" ,
594=> "0001000000000000" ,
595=> "0001000000000000" ,
596=> "0001000000000000" ,
597=> "0001000000000000" ,
598=> "0001000000000000" ,
599=> "0001000000000000" ,
600=> "0001000000000000" ,
601=> "0001000000000000" ,
602=> "0001000000000000" ,
603=> "0001000000000000" ,
604=> "0001000000000000" ,
605=> "0001000000000000" ,
606=> "0001000000000000" ,
607=> "0001000000000000" ,
608=> "0001000000000000" ,
609=> "0001000000000000" ,
610=> "0001000000000000" ,
611=> "0001000000000000" ,
612=> "0001000000000000" ,
613=> "0001000000000000" ,
614=> "0001000000000000" ,
615=> "0001000000000000" ,
616=> "0001000000000000" ,
617=> "0001000000000000" ,
618=> "0001000000000000" ,
619=> "0001000000000000" ,
620=> "0001000000000000" ,
621=> "0001000000000000" ,
622=> "0001000000000000" ,
623=> "0001000000000000" ,
624=> "0001000000000000" ,
625=> "0001000000000000" ,
626=> "0001000000000000" ,
627=> "0001000000000000" ,
628=> "0001000000000000" ,
629=> "0001000000000000" ,
630=> "0001000000000000" ,
631=> "0001000000000000" ,
632=> "0001000000000000" ,
633=> "0001000000000000" ,
634=> "0001000000000000" ,
635=> "0001000000000000" ,
636=> "0001000000000000" ,
637=> "0001000000000000" ,
638=> "0001000000000000" ,
639=> "0001000000000000" ,
640=> "0001000000000000" ,
641=> "0001000000000000" ,
642=> "0001000000000000" ,
643=> "0001000000000000" ,
644=> "0001000000000000" ,
645=> "0001000000000000" ,
646=> "0001000000000000" ,
647=> "0001000000000000" ,
648=> "0001000000000000" ,
649=> "0001000000000000" ,
650=> "0001000000000000" ,
651=> "0001000000000000" ,
652=> "0001000000000000" ,
653=> "0001000000000000" ,
654=> "0001000000000000" ,
655=> "0001000000000000" ,
656=> "0001000000000000" ,
657=> "0001000000000000" ,
658=> "0001000000000000" ,
659=> "0001000000000000" ,
660=> "0001000000000000" ,
661=> "0001000000000000" ,
662=> "0001000000000000" ,
663=> "0001000000000000" ,
664=> "0001000000000000" ,
665=> "0001000000000000" ,
666=> "0001000000000000" ,
667=> "0001000000000000" ,
668=> "0001000000000000" ,
669=> "0001000000000000" ,
670=> "0001000000000000" ,
671=> "0001000000000000" ,
672=> "0001000000000000" ,
673=> "0001000000000000" ,
674=> "0001000000000000" ,
675=> "0001000000000000" ,
676=> "0001000000000000" ,
677=> "0001000000000000" ,
678=> "0001000000000000" ,
679=> "0001000000000000" ,
680=> "0001000000000000" ,
681=> "0001000000000000" ,
682=> "0001000000000000" ,
683=> "0001000000000000" ,
684=> "0001000000000000" ,
685=> "0001000000000000" ,
686=> "0001000000000000" ,
687=> "0001000000000000" ,
688=> "0001000000000000" ,
689=> "0001000000000000" ,
690=> "0001000000000000" ,
691=> "0001000000000000" ,
692=> "0001000000000000" ,
693=> "0001000000000000" ,
694=> "0001000000000000" ,
695=> "0001000000000000" ,
696=> "0001000000000000" ,
697=> "0001000000000000" ,
698=> "0001000000000000" ,
699=> "0001000000000000" ,
700=> "0001000000000000" ,
701=> "0001000000000000" ,
702=> "0001000000000000" ,
703=> "0001000000000000" ,
704=> "0001000000000000" ,
705=> "0001000000000000" ,
706=> "0001000000000000" ,
707=> "0001000000000000" ,
708=> "0001000000000000" ,
709=> "0001000000000000" ,
710=> "0001000000000000" ,
711=> "0001000000000000" ,
712=> "0001000000000000" ,
713=> "0001000000000000" ,
714=> "0001000000000000" ,
715=> "0001000000000000" ,
716=> "0001000000000000" ,
717=> "0001000000000000" ,
718=> "0001000000000000" ,
719=> "0001000000000000" ,
720=> "0001000000000000" ,
721=> "0001000000000000" ,
722=> "0001000000000000" ,
723=> "0001000000000000" ,
724=> "0001000000000000" ,
725=> "0001000000000000" ,
726=> "0001000000000000" ,
727=> "0001000000000000" ,
728=> "0001000000000000" ,
729=> "0001000000000000" ,
730=> "0001000000000000" ,
731=> "0001000000000000" ,
732=> "0001000000000000" ,
733=> "0001000000000000" ,
734=> "0001000000000000" ,
735=> "0001000000000000" ,
736=> "0001000000000000" ,
737=> "0001000000000000" ,
738=> "0001000000000000" ,
739=> "0001000000000000" ,
740=> "0001000000000000" ,
741=> "0001000000000000" ,
742=> "0001000000000000" ,
743=> "0001000000000000" ,
744=> "0001000000000000" ,
745=> "0001000000000000" ,
746=> "0001000000000000" ,
747=> "0001000000000000" ,
748=> "0001000000000000" ,
749=> "0001000000000000" ,
750=> "0001000000000000" ,
751=> "0001000000000000" ,
752=> "0001000000000000" ,
753=> "0001000000000000" ,
754=> "0001000000000000" ,
755=> "0001000000000000" ,
756=> "0001000000000000" ,
757=> "0001000000000000" ,
758=> "0001000000000000" ,
759=> "0001000000000000" ,
760=> "0001000000000000" ,
761=> "0001000000000000" ,
762=> "0001000000000000" ,
763=> "0001000000000000" ,
764=> "0001000000000000" ,
765=> "0001000000000000" ,
766=> "0001000000000000" ,
767=> "0001000000000000" ,
768=> "0000001011110110" ,
769=> "0000001001010001" ,
770=> "0010100000000000" ,
771=> "0001010111000111" ,
772=> "0001000000000000" ,
773=> "0001000000000000" ,
774=> "0001000000000000" ,
775=> "0001000000000000" ,
776=> "0001000000000000" ,
777=> "0001000000000000" ,
778=> "0001000000000000" ,
779=> "0001000000000000" ,
780=> "0001000000000000" ,
781=> "0001000000000000" ,
782=> "0001000000000000" ,
783=> "0001000000000000" ,
784=> "0001000000000000" ,
785=> "0001000000000000" ,
786=> "0001000000000000" ,
787=> "0001000000000000" ,
788=> "0001000000000000" ,
789=> "0001000000000000" ,
790=> "0001000000000000" ,
791=> "0001000000000000" ,
792=> "0001000000000000" ,
793=> "0001000000000000" ,
794=> "0001000000000000" ,
795=> "0001000000000000" ,
796=> "0001000000000000" ,
797=> "0001000000000000" ,
798=> "0001000000000000" ,
799=> "0001000000000000" ,
800=> "0001000000000000" ,
801=> "0001000000000000" ,
802=> "0001000000000000" ,
803=> "0001000000000000" ,
804=> "0001000000000000" ,
805=> "0001000000000000" ,
806=> "0001000000000000" ,
807=> "0001000000000000" ,
808=> "0001000000000000" ,
809=> "0001000000000000" ,
810=> "0001000000000000" ,
811=> "0001000000000000" ,
812=> "0001000000000000" ,
813=> "0001000000000000" ,
814=> "0001000000000000" ,
815=> "0001000000000000" ,
816=> "0001000000000000" ,
817=> "0001000000000000" ,
818=> "0001000000000000" ,
819=> "0001000000000000" ,
820=> "0001000000000000" ,
821=> "0001000000000000" ,
822=> "0001000000000000" ,
823=> "0001000000000000" ,
824=> "0001000000000000" ,
825=> "0001000000000000" ,
826=> "0001000000000000" ,
827=> "0001000000000000" ,
828=> "0001000000000000" ,
829=> "0001000000000000" ,
830=> "0001000000000000" ,
831=> "0001000000000000" ,
832=> "0001000000000000" ,
833=> "0001000000000000" ,
834=> "0001000000000000" ,
835=> "0001000000000000" ,
836=> "0001000000000000" ,
837=> "0001000000000000" ,
838=> "0001000000000000" ,
839=> "0001000000000000" ,
840=> "0001000000000000" ,
841=> "0001000000000000" ,
842=> "0001000000000000" ,
843=> "0001000000000000" ,
844=> "0001000000000000" ,
845=> "0001000000000000" ,
846=> "0001000000000000" ,
847=> "0001000000000000" ,
848=> "0001000000000000" ,
849=> "0001000000000000" ,
850=> "0001000000000000" ,
851=> "0001000000000000" ,
852=> "0001000000000000" ,
853=> "0001000000000000" ,
854=> "0001000000000000" ,
855=> "0001000000000000" ,
856=> "0001000000000000" ,
857=> "0001000000000000" ,
858=> "0001000000000000" ,
859=> "0001000000000000" ,
860=> "0001000000000000" ,
861=> "0001000000000000" ,
862=> "0001000000000000" ,
863=> "0001000000000000" ,
864=> "0001000000000000" ,
865=> "0001000000000000" ,
866=> "0001000000000000" ,
867=> "0001000000000000" ,
868=> "0001000000000000" ,
869=> "0001000000000000" ,
870=> "0001000000000000" ,
871=> "0001000000000000" ,
872=> "0001000000000000" ,
873=> "0001000000000000" ,
874=> "0001000000000000" ,
875=> "0001000000000000" ,
876=> "0001000000000000" ,
877=> "0001000000000000" ,
878=> "0001000000000000" ,
879=> "0001000000000000" ,
880=> "0001000000000000" ,
881=> "0001000000000000" ,
882=> "0001000000000000" ,
883=> "0001000000000000" ,
884=> "0001000000000000" ,
885=> "0001000000000000" ,
886=> "0001000000000000" ,
887=> "0001000000000000" ,
888=> "0001000000000000" ,
889=> "0001000000000000" ,
890=> "0001000000000000" ,
891=> "0001000000000000" ,
892=> "0001000000000000" ,
893=> "0001000000000000" ,
894=> "0001000000000000" ,
895=> "0001000000000000" ,
896=> "0001000000000000" ,
897=> "0001000000000000" ,
898=> "0001000000000000" ,
899=> "0001000000000000" ,
900=> "0001000000000000" ,
901=> "0001000000000000" ,
902=> "0001000000000000" ,
903=> "0001000000000000" ,
904=> "0001000000000000" ,
905=> "0001000000000000" ,
906=> "0001000000000000" ,
907=> "0001000000000000" ,
908=> "0001000000000000" ,
909=> "0001000000000000" ,
910=> "0001000000000000" ,
911=> "0001000000000000" ,
912=> "0001000000000000" ,
913=> "0001000000000000" ,
914=> "0001000000000000" ,
915=> "0001000000000000" ,
916=> "0001000000000000" ,
917=> "0001000000000000" ,
918=> "0001000000000000" ,
919=> "0001000000000000" ,
920=> "0001000000000000" ,
921=> "0001000000000000" ,
922=> "0001000000000000" ,
923=> "0001000000000000" ,
924=> "0001000000000000" ,
925=> "0001000000000000" ,
926=> "0001000000000000" ,
927=> "0001000000000000" ,
928=> "0001000000000000" ,
929=> "0001000000000000" ,
930=> "0001000000000000" ,
931=> "0001000000000000" ,
932=> "0001000000000000" ,
933=> "0001000000000000" ,
934=> "0001000000000000" ,
935=> "0001000000000000" ,
936=> "0001000000000000" ,
937=> "0001000000000000" ,
938=> "0001000000000000" ,
939=> "0001000000000000" ,
940=> "0001000000000000" ,
941=> "0001000000000000" ,
942=> "0001000000000000" ,
943=> "0001000000000000" ,
944=> "0001000000000000" ,
945=> "0001000000000000" ,
946=> "0001000000000000" ,
947=> "0001000000000000" ,
948=> "0001000000000000" ,
949=> "0001000000000000" ,
950=> "0001000000000000" ,
951=> "0001000000000000" ,
952=> "0001000000000000" ,
953=> "0001000000000000" ,
954=> "0001000000000000" ,
955=> "0001000000000000" ,
956=> "0001000000000000" ,
957=> "0001000000000000" ,
958=> "0001000000000000" ,
959=> "0001000000000000" ,
960=> "0001000000000000" ,
961=> "0001000000000000" ,
962=> "0001000000000000" ,
963=> "0001000000000000" ,
964=> "0001000000000000" ,
965=> "0001000000000000" ,
966=> "0001000000000000" ,
967=> "0001000000000000" ,
968=> "0001000000000000" ,
969=> "0001000000000000" ,
970=> "0001000000000000" ,
971=> "0001000000000000" ,
972=> "0001000000000000" ,
973=> "0001000000000000" ,
974=> "0001000000000000" ,
975=> "0001000000000000" ,
976=> "0001000000000000" ,
977=> "0001000000000000" ,
978=> "0001000000000000" ,
979=> "0001000000000000" ,
980=> "0001000000000000" ,
981=> "0001000000000000" ,
982=> "0001000000000000" ,
983=> "0001000000000000" ,
984=> "0001000000000000" ,
985=> "0001000000000000" ,
986=> "0001000000000000" ,
987=> "0001000000000000" ,
988=> "0001000000000000" ,
989=> "0001000000000000" ,
990=> "0001000000000000" ,
991=> "0001000000000000" ,
992=> "0001000000000000" ,
993=> "0001000000000000" ,
994=> "0001000000000000" ,
995=> "0001000000000000" ,
996=> "0001000000000000" ,
997=> "0001000000000000" ,
998=> "0001000000000000" ,
999=> "0001000000000000" ,
1000=> "0001000000000000" ,
1001=> "0001000000000000" ,
1002=> "0001000000000000" ,
1003=> "0001000000000000" ,
1004=> "0001000000000000" ,
1005=> "0001000000000000" ,
1006=> "0001000000000000" ,
1007=> "0001000000000000" ,
1008=> "0001000000000000" ,
1009=> "0001000000000000" ,
1010=> "0001000000000000" ,
1011=> "0001000000000000" ,
1012=> "0001000000000000" ,
1013=> "0001000000000000" ,
1014=> "0001000000000000" ,
1015=> "0001000000000000" ,
1016=> "0001000000000000" ,
1017=> "0001000000000000" ,
1018=> "0001000000000000" ,
1019=> "0001000000000000" ,
1020=> "0001000000000000" ,
1021=> "0001000000000000" ,
1022=> "0001000000000000" ,
1023=> "0001000000000000" ,
1024=> "0001000000000000" ,
1025=> "0001000000000000" ,
1026=> "0001000000000000" ,
1027=> "0001000000000000" ,
1028=> "0001000000000000" ,
1029=> "0001000000000000" ,
1030=> "0001000000000000" ,
1031=> "0001000000000000" ,
1032=> "0001000000000000" ,
1033=> "0001000000000000" ,
1034=> "0001000000000000" ,
1035=> "0001000000000000" ,
1036=> "0001000000000000" ,
1037=> "0001000000000000" ,
1038=> "0001000000000000" ,
1039=> "0001000000000000" ,
1040=> "0001000000000000" ,
1041=> "0001000000000000" ,
1042=> "0001000000000000" ,
1043=> "0001000000000000" ,
1044=> "0001000000000000" ,
1045=> "0001000000000000" ,
1046=> "0001000000000000" ,
1047=> "0001000000000000" ,
1048=> "0001000000000000" ,
1049=> "0001000000000000" ,
1050=> "0001000000000000" ,
1051=> "0001000000000000" ,
1052=> "0001000000000000" ,
1053=> "0001000000000000" ,
1054=> "0001000000000000" ,
1055=> "0001000000000000" ,
1056=> "0001000000000000" ,
1057=> "0001000000000000" ,
1058=> "0001000000000000" ,
1059=> "0001000000000000" ,
1060=> "0001000000000000" ,
1061=> "0001000000000000" ,
1062=> "0001000000000000" ,
1063=> "0001000000000000" ,
1064=> "0001000000000000" ,
1065=> "0001000000000000" ,
1066=> "0001000000000000" ,
1067=> "0001000000000000" ,
1068=> "0001000000000000" ,
1069=> "0001000000000000" ,
1070=> "0001000000000000" ,
1071=> "0001000000000000" ,
1072=> "0001000000000000" ,
1073=> "0001000000000000" ,
1074=> "0001000000000000" ,
1075=> "0001000000000000" ,
1076=> "0001000000000000" ,
1077=> "0001000000000000" ,
1078=> "0001000000000000" ,
1079=> "0001000000000000" ,
1080=> "0001000000000000" ,
1081=> "0001000000000000" ,
1082=> "0001000000000000" ,
1083=> "0001000000000000" ,
1084=> "0001000000000000" ,
1085=> "0001000000000000" ,
1086=> "0001000000000000" ,
1087=> "0001000000000000" ,
1088=> "0001000000000000" ,
1089=> "0001000000000000" ,
1090=> "0001000000000000" ,
1091=> "0001000000000000" ,
1092=> "0001000000000000" ,
1093=> "0001000000000000" ,
1094=> "0001000000000000" ,
1095=> "0001000000000000" ,
1096=> "0001000000000000" ,
1097=> "0001000000000000" ,
1098=> "0001000000000000" ,
1099=> "0001000000000000" ,
1100=> "0001000000000000" ,
1101=> "0001000000000000" ,
1102=> "0001000000000000" ,
1103=> "0001000000000000" ,
1104=> "0001000000000000" ,
1105=> "0001000000000000" ,
1106=> "0001000000000000" ,
1107=> "0001000000000000" ,
1108=> "0001000000000000" ,
1109=> "0001000000000000" ,
1110=> "0001000000000000" ,
1111=> "0001000000000000" ,
1112=> "0001000000000000" ,
1113=> "0001000000000000" ,
1114=> "0001000000000000" ,
1115=> "0001000000000000" ,
1116=> "0001000000000000" ,
1117=> "0001000000000000" ,
1118=> "0001000000000000" ,
1119=> "0001000000000000" ,
1120=> "0001000000000000" ,
1121=> "0001000000000000" ,
1122=> "0001000000000000" ,
1123=> "0001000000000000" ,
1124=> "0001000000000000" ,
1125=> "0001000000000000" ,
1126=> "0001000000000000" ,
1127=> "0001000000000000" ,
1128=> "0001000000000000" ,
1129=> "0001000000000000" ,
1130=> "0001000000000000" ,
1131=> "0001000000000000" ,
1132=> "0001000000000000" ,
1133=> "0001000000000000" ,
1134=> "0001000000000000" ,
1135=> "0001000000000000" ,
1136=> "0001000000000000" ,
1137=> "0001000000000000" ,
1138=> "0001000000000000" ,
1139=> "0001000000000000" ,
1140=> "0001000000000000" ,
1141=> "0001000000000000" ,
1142=> "0001000000000000" ,
1143=> "0001000000000000" ,
1144=> "0001000000000000" ,
1145=> "0001000000000000" ,
1146=> "0001000000000000" ,
1147=> "0001000000000000" ,
1148=> "0001000000000000" ,
1149=> "0001000000000000" ,
1150=> "0001000000000000" ,
1151=> "0001000000000000" ,
1152=> "0001000000000000" ,
1153=> "0001000000000000" ,
1154=> "0001000000000000" ,
1155=> "0001000000000000" ,
1156=> "0001000000000000" ,
1157=> "0001000000000000" ,
1158=> "0001000000000000" ,
1159=> "0001000000000000" ,
1160=> "0001000000000000" ,
1161=> "0001000000000000" ,
1162=> "0001000000000000" ,
1163=> "0001000000000000" ,
1164=> "0001000000000000" ,
1165=> "0001000000000000" ,
1166=> "0001000000000000" ,
1167=> "0001000000000000" ,
1168=> "0001000000000000" ,
1169=> "0001000000000000" ,
1170=> "0001000000000000" ,
1171=> "0001000000000000" ,
1172=> "0001000000000000" ,
1173=> "0001000000000000" ,
1174=> "0001000000000000" ,
1175=> "0001000000000000" ,
1176=> "0001000000000000" ,
1177=> "0001000000000000" ,
1178=> "0001000000000000" ,
1179=> "0001000000000000" ,
1180=> "0001000000000000" ,
1181=> "0001000000000000" ,
1182=> "0001000000000000" ,
1183=> "0001000000000000" ,
1184=> "0001000000000000" ,
1185=> "0001000000000000" ,
1186=> "0001000000000000" ,
1187=> "0001000000000000" ,
1188=> "0001000000000000" ,
1189=> "0001000000000000" ,
1190=> "0001000000000000" ,
1191=> "0001000000000000" ,
1192=> "0001000000000000" ,
1193=> "0001000000000000" ,
1194=> "0001000000000000" ,
1195=> "0001000000000000" ,
1196=> "0001000000000000" ,
1197=> "0001000000000000" ,
1198=> "0001000000000000" ,
1199=> "0001000000000000" ,
1200=> "0001000000000000" ,
1201=> "0001000000000000" ,
1202=> "0001000000000000" ,
1203=> "0001000000000000" ,
1204=> "0001000000000000" ,
1205=> "0001000000000000" ,
1206=> "0001000000000000" ,
1207=> "0001000000000000" ,
1208=> "0001000000000000" ,
1209=> "0001000000000000" ,
1210=> "0001000000000000" ,
1211=> "0001000000000000" ,
1212=> "0001000000000000" ,
1213=> "0001000000000000" ,
1214=> "0001000000000000" ,
1215=> "0001000000000000" ,
1216=> "0001000000000000" ,
1217=> "0001000000000000" ,
1218=> "0001000000000000" ,
1219=> "0001000000000000" ,
1220=> "0001000000000000" ,
1221=> "0001000000000000" ,
1222=> "0001000000000000" ,
1223=> "0001000000000000" ,
1224=> "0001000000000000" ,
1225=> "0001000000000000" ,
1226=> "0001000000000000" ,
1227=> "0001000000000000" ,
1228=> "0001000000000000" ,
1229=> "0001000000000000" ,
1230=> "0001000000000000" ,
1231=> "0001000000000000" ,
1232=> "0001000000000000" ,
1233=> "0001000000000000" ,
1234=> "0001000000000000" ,
1235=> "0001000000000000" ,
1236=> "0001000000000000" ,
1237=> "0001000000000000" ,
1238=> "0001000000000000" ,
1239=> "0001000000000000" ,
1240=> "0001000000000000" ,
1241=> "0001000000000000" ,
1242=> "0001000000000000" ,
1243=> "0001000000000000" ,
1244=> "0001000000000000" ,
1245=> "0001000000000000" ,
1246=> "0001000000000000" ,
1247=> "0001000000000000" ,
1248=> "0001000000000000" ,
1249=> "0001000000000000" ,
1250=> "0001000000000000" ,
1251=> "0001000000000000" ,
1252=> "0001000000000000" ,
1253=> "0001000000000000" ,
1254=> "0001000000000000" ,
1255=> "0001000000000000" ,
1256=> "0001000000000000" ,
1257=> "0001000000000000" ,
1258=> "0001000000000000" ,
1259=> "0001000000000000" ,
1260=> "0001000000000000" ,
1261=> "0001000000000000" ,
1262=> "0001000000000000" ,
1263=> "0001000000000000" ,
1264=> "0001000000000000" ,
1265=> "0001000000000000" ,
1266=> "0001000000000000" ,
1267=> "0001000000000000" ,
1268=> "0001000000000000" ,
1269=> "0001000000000000" ,
1270=> "0001000000000000" ,
1271=> "0001000000000000" ,
1272=> "0001000000000000" ,
1273=> "0001000000000000" ,
1274=> "0001000000000000" ,
1275=> "0001000000000000" ,
1276=> "0001000000000000" ,
1277=> "0001000000000000" ,
1278=> "0001000000000000" ,
1279=> "0001000000000000" ,
1280=> "0001000000000000" ,
1281=> "0001000000000000" ,
OTHERS=>X"0000");

Begin
PROCESS(clk) IS
variable offset: Integer;
BEGIN
	offset:= to_integer(unsigned((address)));
	IF falling_edge(clk) THEN
		IF we = '1' THEN 
			L:for I in 0 to 7 loop
			Li:ram(offset+I) <=  datain(I);
			end loop;
		 END IF;
	END IF;
END PROCESS;
process(address, ram)
	variable offset: Integer;
	BEGIN
	offset:= to_integer(unsigned((address)));
	R:for I in 0 to 7 loop
	Ri:dataout(I) <= ram(offset+I);
	end loop;
end process;

END ARCHITECTURE;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use work.myPackages.all;

Entity CacheSystem is
	port(clk, vrst,rst, MR, MW, MWInstr,int: IN std_logic;
	     address, addressInstr, addressInstrWrite: IN std_logic_vector(10 downto 0);
	     datain: IN std_logic_vector(31 downto 0);
	     PredBits: In std_logic_vector(1 downto 0);
	     instrOut: out std_logic_vector(15 downto 0);
	     dataout: OUT std_logic_vector(31 downto 0));
End CacheSystem;

ARCHITECTURE final of CacheSystem is
signal RamToCach, CachToRam: std_logic;
signal RTCblock, CTRblock: block_Cache;
signal addresstoRam: std_logic_vector(10 downto 0);
signal toInstrCach, ignore: std_logic;
begin
cacheMemoryLabel: entity work.Cache_DataMemory port map(clk, MR, MW, RamToCach, CachToRam, rst,int,address(7 downto 0), datain, dataout, RTCblock, CTRblock);
cacheInstrLabel: entity work.Cache_InstructionMemory port map(clk, MWInstr, toInstrCach, ignore, addressInstr(7 downto 0),addressInstrWrite(7 downto 0),PredBits, instrOut,RTCblock);
cacheControllerLabel: entity work.Cache_Controller port map(clk, vrst,rst, MR, MW, MWInstr, int,address(10 downto 3), addressInstr(10 downto 3), addressInstrwrite(10 downto 3) ,addresstoRam, CachToRam, RamToCach,toInstrCach,ignore);
MainMemoryLabel: entity work.MainMemory port map(clk, CachToRam, addresstoRam, CTRblock, RTCblock);
end ARCHITECTURE;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
 entity test is
	port(clk, rst, MR, MW: IN std_logic;
	     address: IN std_logic_vector(10 downto 0);
	     datain: IN std_logic_vector(31 downto 0);
	     dataout : OUT std_logic_vector(31 downto 0));
End test;

ARCHITECTURE tt of test is
begin
--weeee: entity work.CacheSystem port map(clk, rst, MR, MW, address, datain, dataout);
end tt;

	     